library verilog;
use verilog.vl_types.all;
entity Distributeur_Cafe_vlg_vec_tst is
end Distributeur_Cafe_vlg_vec_tst;
